// nexysA7fpga.sv - Top level module for the Nexys A7 version of the ECE 544 Getting Started project
//
// Created By:	Roy Kravitz
// Date:		26-March-2022
// Version:		2.0
//
// Description:
// ------------
// This module provides the top level for the Getting Started hardware which
// includes the Nexys A7 and no Pmods. Project #1 will add a PmodOLEDrgb and a
// a PmodENC to the system but we didn't want to hold up you working on this
// project while waiting for your Pmods to arrive.
//////////////////////////////////////////////////////////////////////
module nexysA7fpga(
    input logic         clk,			// 100Mhz clock input
    input logic         btnC,			// center pushbutton
    input logic         btnU,			// UP (North) pusbhbutton
    input logic         btnL,			// LEFT (West) pushbutton
    input logic         btnD,			// DOWN (South) pushbutton  - used for system reset
    input logic         btnR,			// RIGHT (East) pushbutton
	input logic         btnCpuReset,	// CPU reset pushbutton
	input logic         encA_0,         // PMOD Encoder A
	input logic         encB_0,         // PMOD Encoder B
	input logic         encBTN_0,       // PMOD Encoder pushbutton
	input logic         encSWT_0,       // PMOD Encoder Switch
    input logic [15:0]  sw,				// slide switches on Nexys 4
    output logic [15:0] led,			// LEDs on Nexys 4   
    output logic        RGB1_Blue,      // RGB1 LED (LD16) 
    output logic        RGB1_Green,
    output logic        RGB1_Red,
    output logic        RGB2_Blue,      // RGB2 LED (LD17)
    output logic        RGB2_Green,
    output logic        RGB2_Red,
    output logic [7:0]  an,             // Seven Segment display
    output logic [6:0]  seg,
    output logic        dp,             // decimal point display on the seven segment 
    
    input logic         uart_rtl_rxd,	// USB UART Rx and Tx on Nexys 4
    output logic        uart_rtl_txd,	
    
	inout logic [3:0]  ja_in,              // JA Pmod 1-4, Inputs from relay (if necessary)
	inout logic [3:0]  ja_out,             // JA Pmod 7-10 Outputs to relay
	inout logic [7:0]  OLED,               // JB Pmod conector - Connected to the PMOD_OLED
	inout logic [3:0]  joystick,           // JC Pmod 1-4, joystick
	inout logic [3:0]  z_step,             // JC Pmod 7-10, Z Stepper
	inout logic [3:0]  x_step,             // JD Pmod 1-4, X Stepper
	inout logic [3:0]  y_step              // JD Pmod 7-10, Y Stepper
	
);

// internal variables
// Clock and Reset 
logic           sysclk; 
logic           sysreset_n, sysreset;

// Joystick pins
logic 		    pmodjstk1_i, pmodjstk1_io, pmodjstk1_o, pmodjstk1_t;
logic 			pmodjstk2_i, pmodjstk2_io, pmodjstk2_o, pmodjstk2_t;
logic 			pmodjstk3_i, pmodjstk3_io, pmodjstk3_o, pmodjstk3_t;
logic 			pmodjstk4_i, pmodjstk4_io, pmodjstk4_o, pmodjstk4_t;

// GPIO Pins
logic [15:0]    gpio_led_out;
logic [4:0]     gpio_btn;
logic [15:0]    gpio_sw;

logic [3:0]    gpio_x_count;
logic [3:0]    gpio_y_count;
logic [3:0]    gpio_z_count;

logic [15:0]    x_cw_cnt;
logic [15:0]    x_ccw_cnt;
logic [15:0]    y_cw_cnt;
logic [15:0]    y_ccw_cnt;
logic [15:0]    z_cw_cnt;
logic [15:0]    z_ccw_cnt;

// OLED pins 
logic 			pmodoledrgb_out_pin1_i, pmodoledrgb_out_pin1_io, pmodoledrgb_out_pin1_o, pmodoledrgb_out_pin1_t; 
logic 			pmodoledrgb_out_pin2_i, pmodoledrgb_out_pin2_io, pmodoledrgb_out_pin2_o, pmodoledrgb_out_pin2_t; 
logic 			pmodoledrgb_out_pin3_i, pmodoledrgb_out_pin3_io, pmodoledrgb_out_pin3_o, pmodoledrgb_out_pin3_t; 
logic 			pmodoledrgb_out_pin4_i, pmodoledrgb_out_pin4_io, pmodoledrgb_out_pin4_o, pmodoledrgb_out_pin4_t; 
logic 			pmodoledrgb_out_pin7_i, pmodoledrgb_out_pin7_io, pmodoledrgb_out_pin7_o, pmodoledrgb_out_pin7_t; 
logic 			pmodoledrgb_out_pin8_i, pmodoledrgb_out_pin8_io, pmodoledrgb_out_pin8_o, pmodoledrgb_out_pin8_t; 
logic 			pmodoledrgb_out_pin9_i, pmodoledrgb_out_pin9_io, pmodoledrgb_out_pin9_o, pmodoledrgb_out_pin9_t; 
logic 			pmodoledrgb_out_pin10_i, pmodoledrgb_out_pin10_io, pmodoledrgb_out_pin10_o, pmodoledrgb_out_pin10_t;

// LED pins 
logic [15:0]    led_int;                // Nexys4IO drives these outputs

// make the connections to the GPIO port.  Most of the bits are unused in the Getting
// Started project but GPIO's provide a convenient way to get the inputs and
// outputs from logic you create to and from the Microblaze.  For example,
// you may decide that using an axi_gpio peripheral is a good way to interface
// your hardware pulse-width detect logic with the Microblaze.  Our application
// is simple.

// Drive the leds from the signal generated by the microblaze 
assign led = led_int;                   // LEDs are driven by led
assign gpio_btn = {encA_0,encB_0,btnC, btnU, btnD, btnL, btnR};
assign gpio_sw = sw;

assign gpio_x_count = x_step;
assign gpio_y_count = y_step;
assign gpio_z_count = z_step;

// make the connections
// system-wide signals
assign sysclk = clk;
assign sysreset_n = btnCpuReset;		// The CPU reset pushbutton is asserted low.  The other pushbuttons are asserted high
										// but the Microblaze for Nexys 4 expects reset to be asserted low
assign sysreset = ~sysreset_n;			// Generate a reset signal that is asserted high for any logic blocks expecting it.

// Pmod OLED connections 
assign OLED[0] = pmodoledrgb_out_pin1_io;
assign OLED[1] = pmodoledrgb_out_pin2_io;
assign OLED[2] = pmodoledrgb_out_pin3_io;
assign OLED[3] = pmodoledrgb_out_pin4_io;
assign OLED[4] = pmodoledrgb_out_pin7_io;
assign OLED[5] = pmodoledrgb_out_pin8_io;
assign OLED[6] = pmodoledrgb_out_pin9_io;
assign OLED[7] = pmodoledrgb_out_pin10_io;

// JA can be used for debug purposes
//assign JA = 8'b0000000;

// Pmodjstk2 signals
// JC - top row
assign  pmodjstk1_io = joystick[0];
assign  pmodjstk2_io = joystick[1];
assign  pmodjstk3_io = joystick[2];
assign  pmodjstk4_io = joystick[3];

// instantiate the embedded system
embsys EMBSYS
(
        // RGB1/2 Led's 
        .RGB1_Blue_0(RGB1_Blue),
        .RGB1_Green_0(RGB1_Green),
        .RGB1_Red_0(RGB1_Red),
        .RGB2_Blue_0(RGB2_Blue),
        .RGB2_Green_0(RGB2_Green),
        .RGB2_Red_0(RGB2_Red),
        
         // Seven Segment Display anode control  
        .an_0(an),
        .dp_0(dp),
        //.led_0(led_int),
        .seg_0(seg),

        // PMOD JSTCK
        .jc_1_4_pin1_i(pmodjstk1_i),
        .jc_1_4_pin1_o(pmodjstk1_o),
        .jc_1_4_pin1_t(pmodjstk1_t),
        .jc_1_4_pin2_i(pmodjstk2_i),
        .jc_1_4_pin2_o(pmodjstk2_o),
        .jc_1_4_pin2_t(pmodjstk2_t),
        .jc_1_4_pin3_i(pmodjstk3_i),
        .jc_1_4_pin3_o(pmodjstk3_o),
        .jc_1_4_pin3_t(pmodjstk3_t),
        .jc_1_4_pin4_i(pmodjstk4_i),
        .jc_1_4_pin4_o(pmodjstk4_o),
        .jc_1_4_pin4_t(pmodjstk4_t),
        
        // PMOD OLED pins 
        .jb_pin10_i(pmodoledrgb_out_pin10_i),
	    .jb_pin10_o(pmodoledrgb_out_pin10_o),
	    .jb_pin10_t(pmodoledrgb_out_pin10_t),
	    .jb_pin1_i(pmodoledrgb_out_pin1_i),
	    .jb_pin1_o(pmodoledrgb_out_pin1_o),
	    .jb_pin1_t(pmodoledrgb_out_pin1_t),
	    .jb_pin2_i(pmodoledrgb_out_pin2_i),
	    .jb_pin2_o(pmodoledrgb_out_pin2_o),
	    .jb_pin2_t(pmodoledrgb_out_pin2_t),
	    .jb_pin3_i(pmodoledrgb_out_pin3_i),
	    .jb_pin3_o(pmodoledrgb_out_pin3_o),
	    .jb_pin3_t(pmodoledrgb_out_pin3_t),
	    .jb_pin4_i(pmodoledrgb_out_pin4_i),
	    .jb_pin4_o(pmodoledrgb_out_pin4_o),
	    .jb_pin4_t(pmodoledrgb_out_pin4_t),
	    .jb_pin7_i(pmodoledrgb_out_pin7_i),
	    .jb_pin7_o(pmodoledrgb_out_pin7_o),
	    .jb_pin7_t(pmodoledrgb_out_pin7_t),
	    .jb_pin8_i(pmodoledrgb_out_pin8_i),
	    .jb_pin8_o(pmodoledrgb_out_pin8_o),
	    .jb_pin8_t(pmodoledrgb_out_pin8_t),
	    .jb_pin9_i(pmodoledrgb_out_pin9_i),
	    .jb_pin9_o(pmodoledrgb_out_pin9_o),
	    .jb_pin9_t(pmodoledrgb_out_pin9_t),
	    
	    // GPIO Inputs and Outputs
	    .gpio_led_tri_o(led_int),
	    .gpio_btn_tri_i(gpio_btn),
        .gpio_sw_tri_i(gpio_sw),
        
        // GPIO for counting X, Y, and Z
        .x_count_tri_i(gpio_x_count),
        .y_count_tri_i(gpio_y_count),
        .z_count_tri_i(gpio_z_count),
       
        //JA Inputs/Outputs
        .gpio_ja_1_4_in_tri_i(ja_in),
        .gpio_ja_7_10_out_tri_o(ja_out),
        
        // X Count Outputs
        .x_cw_cnt_0(x_cw_cnt),
        .x_ccw_cnt_0(x_ccw_cnt),
        
        // Y Count Outputs
        .y_cw_cnt_0(y_cw_cnt),
        .y_ccw_cnt_0(y_ccw_cnt),
        
        // Z Count Outputs
        .z_cw_cnt_0(z_cw_cnt),
        .z_ccw_cnt_0(z_ccw_cnt),
        
        // Stepper Outputs
        .jc_7_10(z_step),
        .jd_1_4(x_step),
        .jd_7_10(y_step),
        
        // Push buttons and switches  
        .btnC_0(btnC),
        .btnD_0(btnD),
        .btnL_0(btnL),
        .btnR_0(btnR),
        .btnU_0(btnU),
        .sw_0(sw),
        
        // reset and clock 
        .sysreset_n(sysreset_n),
        .sysclk(sysclk),
        
        // UART pins 
        .usb_uart_rxd(uart_rtl_rxd),
        .usb_uart_txd(uart_rtl_txd)
);
 
// Tristate buffers for the pmodOLEDrgb pins
// generated by PMOD bridge component.  Many
// of these signals are not tri-state.
IOBUF pmodoledrgb_out_pin1_iobuf
(
    .I(pmodoledrgb_out_pin1_o),
    .IO(pmodoledrgb_out_pin1_io),
    .O(pmodoledrgb_out_pin1_i),
    .T(pmodoledrgb_out_pin1_t)
);

IOBUF pmodoledrgb_out_pin2_iobuf
(
    .I(pmodoledrgb_out_pin2_o),
    .IO(pmodoledrgb_out_pin2_io),
    .O(pmodoledrgb_out_pin2_i),
    .T(pmodoledrgb_out_pin2_t)
);

IOBUF pmodoledrgb_out_pin3_iobuf
(
    .I(pmodoledrgb_out_pin3_o),
    .IO(pmodoledrgb_out_pin3_io),
    .O(pmodoledrgb_out_pin3_i),
    .T(pmodoledrgb_out_pin3_t)
);

IOBUF pmodoledrgb_out_pin4_iobuf
(
    .I(pmodoledrgb_out_pin4_o),
    .IO(pmodoledrgb_out_pin4_io),
    .O(pmodoledrgb_out_pin4_i),
    .T(pmodoledrgb_out_pin4_t)
);

IOBUF pmodoledrgb_out_pin7_iobuf
(
    .I(pmodoledrgb_out_pin7_o),
    .IO(pmodoledrgb_out_pin7_io),
    .O(pmodoledrgb_out_pin7_i),
    .T(pmodoledrgb_out_pin7_t)
);

IOBUF pmodoledrgb_out_pin8_iobuf
(
    .I(pmodoledrgb_out_pin8_o),
    .IO(pmodoledrgb_out_pin8_io),
    .O(pmodoledrgb_out_pin8_i),
    .T(pmodoledrgb_out_pin8_t)
);

IOBUF pmodoledrgb_out_pin9_iobuf
(
    .I(pmodoledrgb_out_pin9_o),
    .IO(pmodoledrgb_out_pin9_io),
    .O(pmodoledrgb_out_pin9_i),
    .T(pmodoledrgb_out_pin9_t)
);

IOBUF pmodoledrgb_out_pin10_iobuf
(
    .I(pmodoledrgb_out_pin10_o),
    .IO(pmodoledrgb_out_pin10_io),
    .O(pmodoledrgb_out_pin10_i),
    .T(pmodoledrgb_out_pin10_t)
);

// Tristate buffers for the pmodCompass pins
// generated by PMOD bridge component.  Many
// of these signals are not tri-state.
IOBUF pmodjstk1_iobuf
     (.I(pmodjstk1_o),
      .IO(pmodjstk1_io),
      .O(pmodjstk1_i),
      .T(pmodjstk1_t));
	  
IOBUF pmodjstk2_iobuf
     (.I(pmodjstk2_o),
      .IO(pmodjstk2_io),
      .O(pmodjstk2_i),
      .T(pmodjstk2_t));
	  
IOBUF pmodjstk3_iobuf
     (.I(pmodjstk3_o),
      .IO(pmodjstk3_io),
      .O(pmodjstk3_i),
      .T(pmodjstk3_t));
	  
IOBUF pmodjstk4_iobuf
     (.I(pmodjstk4_o),
      .IO(pmodjstk4_io),
      .O(pmodjstk4_i),
      .T(pmodjstk4_t));

endmodule: nexysA7fpga


